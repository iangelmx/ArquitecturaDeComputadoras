
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity PROCESADOR_ESCOMIPS is
	Port(
		clk, clr : in STD_LOGIC;
		read_data2 : out STD_LOGIC_VECTOR (15 downto 0)
	);
end PROCESADOR_ESCOMIPS;

architecture Behavioral of PROCESADOR_ESCOMIPS is

begin


end Behavioral;

