
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package ESCOMIPS_lib is



end ESCOMIPS_lib;

package body ESCOMIPS_lib is


 
end ESCOMIPS_lib;
